// PLLClk.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module PLLClk (
		output wire  pll_0_outclk0_clk, // pll_0_outclk0.clk
		input  wire  pll_0_refclk_clk,  //  pll_0_refclk.clk
		input  wire  pll_0_reset_reset  //   pll_0_reset.reset
	);

	PLLClk_pll_0 pll_0 (
		.refclk   (pll_0_refclk_clk),  //  refclk.clk
		.rst      (pll_0_reset_reset), //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.locked   ()                   // (terminated)
	);

endmodule
